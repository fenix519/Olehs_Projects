** Profile: "SCHEMATIC1-PFET charge"  [ O:\SPICE\PFET-Input_Charge_r00\pfet_input_charge-pspicefiles\schematic1\pfet charge.sim ] 

** Creating circuit file "PFET charge.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "O:/SPICE/tpc6130.lib" 
.LIB "D:/Programs/Cadence/SPB_17.2/tools/capture/library/pspice/infineon_optimos_p.olb" 
.LIB "O:/SPICE/ssm6p49nu_pspice_20140521.lib" 
* From [PSPICE NETLIST] section of C:\Users\nazar\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2m 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
